`include "defines.v"


module pipectrl(
    input wire clk_i,
    input wire rs1_i,
    



);




endmodule